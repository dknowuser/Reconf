// nios_tb.v

// Generated using ACDS version 12.1sp1 243 at 2020.10.10.18:17:48

`timescale 1 ps / 1 ps
module nios_tb (
	);

	wire        nios_inst_clk_bfm_clk_clk;                  // nios_inst_clk_bfm:clk -> nios_inst:clk_clk
	wire  [7:0] nios_inst_pio_0_external_connection_export; // nios_inst:pio_0_external_connection_export -> nios_inst_pio_0_external_connection_bfm:sig_export

	nios nios_inst (
		.clk_clk                          (nios_inst_clk_bfm_clk_clk),                  //                       clk.clk
		.pio_0_external_connection_export (nios_inst_pio_0_external_connection_export)  // pio_0_external_connection.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_inst_clk_bfm (
		.clk (nios_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm nios_inst_pio_0_external_connection_bfm (
		.sig_export (nios_inst_pio_0_external_connection_export)  // conduit.export
	);

endmodule
